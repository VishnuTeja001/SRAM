


package s_ram_pkg_file;

`include "uvm_pkg.sv"

import uvm_pkg::*;

	
`include "mem_seq_item.sv"
`include "mem_sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "mem_omonitor.sv"
`include "agent_1.sv"
`include "scoreboard.sv"
//`include  "scbd_2ap.sv"
//`include  "scbd_get_fifo.sv"
`include "environment.sv"
//`include  "env_2ap.sv"
`include "test.sv"


endpackage
